module add4 (
    add4i, add4o
);
input [31:0] add4i;
output [31:0] add4o;

assign add4o = add4i +4;

endmodule